../../../../../../RuflCore/firmware/hdl/ReuseableElements/DataPipe64.vhd