../../../../../../RuflCore/firmware/hdl/ReuseableElements/DataPipe32.vhd