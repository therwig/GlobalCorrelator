../../../../../../RuflCore/firmware/hdl/ReuseableElements/DataPipe128.vhd