../../../../../../RuflCore/firmware/hdl/ReuseableElements/DataPipeN.vhd