../../../../../../RuflCore/firmware/hdl/ReuseableElements/DataPipe16.vhd